localparam FUNCT_ADD_RAW    = 10'b0000000000;
localparam FUNCT_SUB_RAW    = 10'b0100000000;
localparam FUNCT_OR_RAW     = 10'b0000000110;
localparam FUNCT_XOR_RAW    = 10'b0000000100;
localparam FUNCT_AND_RAW    = 10'b0000000111;
localparam FUNCT_SLT_RAW    = 10'b0000000010;
localparam FUNCT_SLTU_RAW   = 10'b0000000011;
localparam FUNCT_SLL_RAW    = 10'b0000000001;
localparam FUNCT_SRL_RAW    = 10'b0000000101;
localparam FUNCT_SRA_RAW    = 10'b0100000101;

localparam FUNCT_NOP_OH     = 10'b0000000000;
localparam FUNCT_ADD_OH     = 10'b0000000001;
localparam FUNCT_SUB_OH     = 10'b0000000010;
localparam FUNCT_OR_OH      = 10'b0000000100;
localparam FUNCT_XOR_OH     = 10'b0000001000;
localparam FUNCT_AND_OH     = 10'b0000010000;
localparam FUNCT_STL_OH     = 10'b0000100000;
localparam FUNCT_STLU_OH    = 10'b0001000000;
localparam FUNCT_SLL_OH     = 10'b0010000000;
localparam FUNCT_SRL_OH     = 10'b0100000000;
localparam FUNCT_SRA_OH     = 10'b1000000000;

localparam MEM_FUNCT_LB_RAW  = 3'b000;
localparam MEM_FUNCT_LH_RAW  = 3'b001;
localparam MEM_FUNCT_LW_RAW  = 3'b010;
localparam MEM_FUNCT_LBU_RAW = 3'b100;
localparam MEM_FUNCT_LHU_RAW = 3'b101;
//Decoded in seperate processes
localparam MEM_FUNCT_SB_RAW  = 3'b000;
localparam MEM_FUNCT_SH_RAW  = 3'b001;
localparam MEM_FUNCT_SW_RAW  = 3'b010;

localparam MEM_FUNCT_NOP_OH = 8'b00000000;
localparam MEM_FUNCT_LB_OH  = 8'b00000001;
localparam MEM_FUNCT_LH_OH  = 8'b00000010;
localparam MEM_FUNCT_LW_OH  = 8'b00000100;
localparam MEM_FUNCT_LBU_OH = 8'b00001000;
localparam MEM_FUNCT_LHU_OH = 8'b00010000;
localparam MEM_FUNCT_SB_OH  = 8'b00100000;
localparam MEM_FUNCT_SH_OH  = 8'b01000000;
localparam MEM_FUNCT_SW_OH  = 8'b10000000;

localparam BR_FUNCT_BEQ_RAW  = 3'b000;
localparam BR_FUNCT_BNE_RAW  = 3'b001;
localparam BR_FUNCT_BLT_RAW  = 3'b100;
localparam BR_FUNCT_BGE_RAW  = 3'b101;
localparam BR_FUNCT_BLTU_RAW = 3'b110;
localparam BR_FUNCT_BGEU_RAW = 3'b111;

localparam BR_FUNCT_NOP_OH  = 7'b0000000;
localparam BR_FUNCT_BEQ_OH  = 7'b0000001;
localparam BR_FUNCT_BNE_OH  = 7'b0000010;
localparam BR_FUNCT_BLT_OH  = 7'b0000100;
localparam BR_FUNCT_BGE_OH  = 7'b0001000;
localparam BR_FUNCT_BLTU_OH = 7'b0010000;
localparam BR_FUNCT_BGEU_OH = 7'b0100000;
//Handles JALR and JAL
localparam BR_FUNCT_JUMP_OH = 7'b1000000;
